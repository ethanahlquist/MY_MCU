`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Bridget Benson 
// 
// Create Date: 10/01/2018 10:22:13 AM
// Description: Generic Clock Divider.  Divides the input clock by MAXCOUNT*2
// 
//////////////////////////////////////////////////////////////////////////////////


module ClockDivider (
    input clk, 
    input [16:0] maxcount,
    output logic sclk = 0
    );     
        
    logic [16:0] count = 0; 
    
    always_ff @ (posedge clk)
    begin
        count = count +2;  // this count is supposed to restart at half the period, so we essentially divide period by two.

        if(maxcount == 0)
        begin
            //count = 0;
            sclk = 0;
        end
        else if (count >= maxcount)
        begin
            count = 0;
            sclk = ~sclk;
        end
             
    end
    
endmodule