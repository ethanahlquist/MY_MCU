`timescale 1ns / 1ps

module MORE_TEMP_TOP(
input BTNR,
input BTNU,
input BTNL,
input BTND,
output logic [4:0] BUTTONS
    );
    
    //temp_top temp_top(.*);
    
    //RAT_MCU MCU(.*);
    //FLAGS FLAGS(.*);
    //STACK_POINTER SP(.*);
    //RAT_WRAPPER TOP(.*);
    
endmodule
